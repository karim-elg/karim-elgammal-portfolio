-- Simple OR gate design

--Import statements of the libraries used
library IEEE;
use IEEE.std_logic_1164.all;


--Decleration of the 'black box' or_gate
entity or_gate is
port(
  a: in std_logic;
  b: in std_logic;
  q: out std_logic);
end or_gate;

--Structural behaviour of the or_gate entity

architecture rtl of or_gate is
begin
  process(a, b) is
  begin
    q <= a or b;
  end process;
end rtl;
